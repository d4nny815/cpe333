

module top;

cam_itf itf();
testbench tb(.*);
grader gdr(.*);

endmodule : top
