import mult_types::*;

module top;
    multiplier_itf itf();
    testbench tb (.*);
    grader grd (.*);
endmodule : top
