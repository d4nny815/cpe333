`timescale 1ns / 1ps

module instr_cache (
    input [31:0] addr_i,
    input [31:0] data_i,
    input reset,
    output hit,
    output [31:0] data_o,
    output [31:0] addr_o,
    output dirty_o
)


endmodule