    Mac OS X            	   2  �     �                                    ATTR���a  �   �   :                  �   :  com.apple.quarantine 0081;6564fb82;Firefox;3FE77678-00C9-43AF-A061-D6AF481826A2                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             This resource fork intentionally left blank                                                                                                                                                                                                                            ��