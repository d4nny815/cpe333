module cacheline_adaptor
(
    mem_itf.device ca_itf,
    mem_itf.controller pmem_itf
);

 

endmodule : cacheline_adaptor